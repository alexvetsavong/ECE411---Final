// Wallace Tree Multiplier