import rv32i_types::*;

module datapath();
// TODO: create control_rom module

// TODO: instantiate modules for each stage

// IF


// ID


// EX


// MEM


// WB


endmodule